`ifndef __RSA_DEFINE__
`define __RSA_DEFINE__

// 128, 256, 512, 1024

parameter RSA_MAX = 1024;
parameter RSA_BUS = (RSA_MAX-1);
parameter RSA_MAX_LOG2 = 12;

//parameter RSA_BIT = 256;
//parameter RSA_CHUNK = RSA_BIT/8;

`endif