`include "include/RecorderDefine.vh"

module OutputController(
    input           i_clk,
    input           i_rst,
    // Recorder Core
    input   [15:0]  i_output_event,
    input   [23:0]  i_time
    // LCD Controller
);

endmodule